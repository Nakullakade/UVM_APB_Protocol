package apb_package;
`include "uvm_macros.svh" 
 import uvm_pkg::*;

`include "apb_sequence_item.sv"
`include "apb_slave_monitor.sv"
`include "apb_master_monitor.sv"
`include "apb_master_driver.sv"
`include "apb_master_sequencer.sv"
`include "master_agent_config.sv"
`include "slave_agent_config.sv"
`include "env_config.sv"
`include "apb_slave_agent.sv"
`include "apb_master_agent.sv"
`include "apb_scoreboard.sv"
`include "apb_functional_coverage.sv"
`include "apb_virtual_sequencer.sv"
`include "apb_environment.sv"
`include "apb_sequence.sv"
`include "apb_virtual_sequence.sv"
`include "apb_test.sv"
endpackage